----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/01/2022 05:40:37 PM
-- Design Name: 
-- Module Name: embedded_kcpsm6 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity embedded_kcpsm6 is
  port (                   
                             in_port : in std_logic_vector(7 downto 0);
                            out_port : out std_logic_vector(7 downto 0);
                             port_id : out std_logic_vector(7 downto 0);
                        write_strobe : out std_logic;
                      --k_write_strobe : out std_logic;
                        -- read_strobe : out std_logic;
                           --interrupt : in std_logic;
                       --interrupt_ack : out std_logic;
                           --    sleep : in std_logic;
                                 clk : in std_logic;
                                 rst : in std_logic);
end embedded_kcpsm6;

architecture Behavioral of embedded_kcpsm6 is

component kcpsm6 
    generic(                 hwbuild : std_logic_vector(7 downto 0) := X"00";
                    interrupt_vector : std_logic_vector(11 downto 0) := X"3FF";
             scratch_pad_memory_size : integer := 64);
    port (                   address : out std_logic_vector(11 downto 0);
                         instruction : in std_logic_vector(17 downto 0);
                         bram_enable : out std_logic;
                             in_port : in std_logic_vector(7 downto 0);
                            out_port : out std_logic_vector(7 downto 0);
                             port_id : out std_logic_vector(7 downto 0);
                        write_strobe : out std_logic;
                      k_write_strobe : out std_logic;
                         read_strobe : out std_logic;
                           interrupt : in std_logic;
                       interrupt_ack : out std_logic;
                               sleep : in std_logic;
                               reset : in std_logic;
                                 clk : in std_logic);
end component;

component your_program is
    Port (      address : in std_logic_vector(11 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                 enable : in std_logic;
                    clk : in std_logic);
end component;

-- Signals for connection of KCPSM6 and Program Memory.
--

signal           address : std_logic_vector(11 downto 0);
signal       instruction : std_logic_vector(17 downto 0);
signal       bram_enable : std_logic;
signal       interrupt_s : std_logic;
signal   interrupt_ack_s : std_logic;
signal      kcpsm6_sleep : std_logic;
signal      kcpsm6_reset : std_logic;

begin


processor: kcpsm6
    generic map (                 hwbuild => X"00", 
                         interrupt_vector => X"3FF",
                  scratch_pad_memory_size => 64)
    port map(      address => address,
               instruction => instruction,
               bram_enable => bram_enable,
                   port_id => port_id,
              write_strobe => write_strobe,
            k_write_strobe => open,
                  out_port => out_port,
               read_strobe => open,
                   in_port => in_port,
                 interrupt => interrupt_s,
             interrupt_ack => interrupt_ack_s,
                     sleep => kcpsm6_sleep,
                     reset => kcpsm6_reset,
                       clk => clk);
                       
program_rom: your_program                    --Name to match your PSM file
 
    port map(      address => address,      
               instruction => instruction,
                    enable => bram_enable,
                       clk => clk);

kcpsm6_reset <= rst;
kcpsm6_sleep <= '0';
interrupt_s <= interrupt_ack_s; 

end Behavioral;
